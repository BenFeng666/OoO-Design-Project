module ALU(
    input wire [31:0] A,
    input wire [31:0] B,
    input wire [3:0] ctrl,
    output reg [31:0] result,
    output reg zero,
    output reg negative

);

always @(*) begin
    case (ctrl)
    4'b0000: result = A+B;
    4'b0001: result = A-B;
    4'b0010: result = A&B;
    4'b0011: result = A|B;
    4'b0100: result = A^B;
    4'b0101: result = A << B[4:0];
    4'b0110: result = A>>B[4:0];
    4'b0111: result = $signed(A)>>>B[4:0];
    4'b1000: result = ($signed(A)<$signed(B))? 32'd1:32'd0;
    4'b1001: result = (A<B)? 32'd1:32'd0;
    default: result=32'b0; 
    endcase

    if (result == 32'b0)begin
      zero=1;
    end
    else begin
        zero=0 ;
    end
    
    negative = result[31]; 


end

endmodule
